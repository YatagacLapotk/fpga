module and_gate (
    input wire in1, in2,
    output wire out1
);

    assign out1 = in1 & in2;
    
endmodule